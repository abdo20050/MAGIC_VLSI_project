magic
tech scmos
timestamp 1667779387
<< metal1 >>
rect -28 20 12 24
rect 56 20 96 24
rect 56 0 60 4
rect -56 -4 -52 0
rect -16 -4 -12 0
<< metal2 >>
rect -56 60 120 64
rect -56 56 -52 60
rect 116 56 120 60
rect -16 52 80 56
rect 0 40 4 44
<< m2contact >>
rect -32 20 -28 24
rect 96 20 100 24
use trans2to1  trans2to1_0
timestamp 1664050318
transform 1 0 4 0 1 0
box -4 0 60 44
use trans2to1  trans2to1_1
timestamp 1664050318
transform 0 1 76 -1 0 52
box -4 0 60 44
use trans2to1  trans2to1_2
timestamp 1664050318
transform 0 -1 -12 -1 0 52
box -4 0 60 44
<< end >>

magic
tech scmos
timestamp 1664037220
<< metal1 >>
rect -20 57 -16 108
rect -8 68 0 72
rect 108 47 112 100
rect -24 32 0 36
rect -60 -19 -48 -15
rect -60 -83 -56 -19
rect -12 -44 -8 0
rect 80 -7 84 43
rect 159 4 168 8
rect 88 -24 91 2
rect 64 -28 91 -24
rect 0 -56 4 -51
rect -8 -60 4 -56
rect -60 -86 0 -83
<< metal2 >>
rect -16 108 8 112
rect 4 104 8 108
rect 72 100 108 104
rect 84 43 95 47
rect 64 20 91 24
rect -8 0 0 4
rect 72 -11 80 -7
rect -16 -47 -12 -44
rect -20 -48 -12 -47
rect -20 -107 -16 -48
rect 95 -107 100 -57
rect -20 -111 0 -107
rect 72 -111 100 -107
<< m2contact >>
rect -20 108 -16 112
rect 108 100 112 104
rect -20 53 -16 57
rect 80 43 84 47
rect 108 43 112 47
rect 60 20 64 24
rect -12 0 -8 4
rect 91 20 95 24
rect 80 -11 84 -7
rect -12 -48 -8 -44
use and  and_0
timestamp 1663595043
transform 1 0 0 0 1 0
box 0 0 72 104
use and  and_1
timestamp 1663595043
transform 1 0 0 0 1 -111
box 0 0 72 104
use not  not_0
timestamp 1663582360
transform 1 0 -56 0 1 -47
box 8 0 40 104
use or  or_0
timestamp 1663598260
transform 1 0 91 0 1 -57
box 0 0 76 104
<< end >>

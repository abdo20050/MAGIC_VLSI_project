magic
tech scmos
timestamp 1667974587
<< polysilicon >>
rect 2366 303 2368 307
rect 2346 301 2348 303
rect 2352 301 2424 303
rect 2428 301 2430 303
rect 2382 288 2384 291
rect 2346 286 2348 288
rect 2352 286 2424 288
rect 2428 286 2430 288
rect 2410 241 2412 249
rect 2342 239 2344 241
rect 2348 239 2428 241
rect 2432 239 2434 241
rect 2357 196 2360 200
rect 2346 194 2348 196
rect 2352 194 2424 196
rect 2428 194 2430 196
rect 2346 182 2348 184
rect 2352 182 2412 184
rect 2416 182 2424 184
rect 2428 182 2430 184
rect 2410 152 2412 160
rect 2342 150 2344 152
rect 2348 150 2428 152
rect 2432 150 2434 152
rect 2410 109 2412 117
rect 2342 107 2344 109
rect 2348 107 2428 109
rect 2432 107 2434 109
rect 2366 68 2368 72
rect 2346 66 2348 68
rect 2352 66 2424 68
rect 2428 66 2430 68
rect 2382 53 2384 56
rect 2346 51 2348 53
rect 2352 51 2424 53
rect 2428 51 2430 53
rect 2410 15 2412 23
rect 2342 13 2344 15
rect 2348 13 2428 15
rect 2432 13 2434 15
rect 2357 -20 2360 -16
rect 2346 -22 2348 -20
rect 2352 -22 2424 -20
rect 2428 -22 2430 -20
rect 2346 -34 2348 -32
rect 2352 -34 2412 -32
rect 2416 -34 2424 -32
rect 2428 -34 2430 -32
rect 2410 -64 2412 -56
rect 2342 -66 2344 -64
rect 2348 -66 2428 -64
rect 2432 -66 2434 -64
rect 2410 -102 2412 -94
rect 2342 -104 2344 -102
rect 2348 -104 2428 -102
rect 2432 -104 2434 -102
rect 2366 -139 2368 -135
rect 2346 -141 2348 -139
rect 2352 -141 2424 -139
rect 2428 -141 2430 -139
rect 2382 -154 2384 -151
rect 2346 -156 2348 -154
rect 2352 -156 2424 -154
rect 2428 -156 2430 -154
<< ndiffusion >>
rect 2424 311 2428 315
rect 2424 303 2428 307
rect 2424 299 2428 301
rect 2424 288 2428 295
rect 2424 283 2428 286
rect 2424 275 2428 279
rect 2428 249 2432 253
rect 2428 241 2432 245
rect 2428 233 2432 239
rect 2428 225 2432 229
rect 2424 196 2428 200
rect 2424 184 2428 194
rect 2424 172 2428 182
rect 2428 160 2432 164
rect 2428 152 2432 156
rect 2428 144 2432 150
rect 2428 136 2432 140
rect 2428 117 2432 121
rect 2428 109 2432 113
rect 2428 101 2432 107
rect 2428 93 2432 97
rect 2424 76 2428 80
rect 2424 68 2428 72
rect 2424 64 2428 66
rect 2424 53 2428 60
rect 2424 48 2428 51
rect 2424 40 2428 44
rect 2428 23 2432 27
rect 2428 15 2432 19
rect 2428 7 2432 13
rect 2428 -1 2432 3
rect 2424 -20 2428 -16
rect 2424 -32 2428 -22
rect 2424 -44 2428 -34
rect 2428 -56 2432 -52
rect 2428 -64 2432 -60
rect 2428 -72 2432 -66
rect 2428 -80 2432 -76
rect 2428 -94 2432 -90
rect 2428 -102 2432 -98
rect 2428 -110 2432 -104
rect 2428 -118 2432 -114
rect 2424 -131 2428 -127
rect 2424 -139 2428 -135
rect 2424 -143 2428 -141
rect 2424 -154 2428 -147
rect 2424 -159 2428 -156
rect 2424 -167 2428 -163
<< pdiffusion >>
rect 2348 311 2352 315
rect 2348 303 2352 307
rect 2348 288 2352 301
rect 2348 283 2352 286
rect 2348 275 2352 279
rect 2344 249 2348 253
rect 2344 241 2348 245
rect 2344 233 2348 239
rect 2344 225 2348 229
rect 2348 196 2352 200
rect 2348 192 2352 194
rect 2348 184 2352 188
rect 2348 176 2352 182
rect 2348 168 2352 172
rect 2344 160 2348 164
rect 2344 152 2348 156
rect 2344 144 2348 150
rect 2344 136 2348 140
rect 2344 117 2348 121
rect 2344 109 2348 113
rect 2344 101 2348 107
rect 2344 93 2348 97
rect 2348 76 2352 80
rect 2348 68 2352 72
rect 2348 53 2352 66
rect 2348 48 2352 51
rect 2348 40 2352 44
rect 2344 23 2348 27
rect 2344 15 2348 19
rect 2344 7 2348 13
rect 2344 -1 2348 3
rect 2348 -20 2352 -16
rect 2348 -24 2352 -22
rect 2348 -32 2352 -28
rect 2348 -40 2352 -34
rect 2348 -48 2352 -44
rect 2344 -56 2348 -52
rect 2344 -64 2348 -60
rect 2344 -72 2348 -66
rect 2344 -80 2348 -76
rect 2344 -94 2348 -90
rect 2344 -102 2348 -98
rect 2344 -110 2348 -104
rect 2344 -118 2348 -114
rect 2348 -131 2352 -127
rect 2348 -139 2352 -135
rect 2348 -154 2352 -141
rect 2348 -159 2352 -156
rect 2348 -167 2352 -163
<< metal1 >>
rect 2248 792 2252 980
rect -892 705 -881 709
rect -892 436 -888 705
rect -848 336 -844 693
rect -704 452 -700 621
rect -412 617 -405 621
rect -400 552 -396 721
rect 615 721 680 725
rect -392 705 -385 709
rect -392 428 -388 705
rect -348 344 -344 689
rect -192 460 -188 621
rect 20 56 24 548
rect 116 544 120 721
rect 140 709 151 713
rect 104 188 108 432
rect 140 420 144 709
rect 128 240 132 284
rect 148 228 152 332
rect 184 196 188 348
rect 192 336 196 697
rect 163 192 188 196
rect 204 136 208 203
rect 156 52 160 132
rect 236 80 240 540
rect 372 468 376 621
rect 676 536 680 721
rect 1656 721 1680 725
rect 692 712 699 716
rect 300 188 304 424
rect 324 240 328 292
rect 344 228 348 340
rect 380 200 384 356
rect 360 196 384 200
rect 396 124 400 203
rect 200 56 204 76
rect 340 52 344 120
rect 432 80 436 532
rect 468 188 472 416
rect 492 240 496 300
rect 512 228 516 332
rect 552 200 556 364
rect 528 196 556 200
rect 564 112 568 203
rect 380 56 384 76
rect 520 52 524 108
rect 592 80 596 524
rect 692 412 696 712
rect 648 188 652 408
rect 732 328 736 697
rect 672 240 676 308
rect 692 228 696 324
rect 740 200 744 372
rect 708 196 744 200
rect 748 100 752 203
rect 560 56 564 76
rect 700 52 704 96
rect 788 84 792 512
rect 896 476 900 621
rect 1192 528 1196 721
rect 1199 712 1203 713
rect 844 188 848 268
rect 868 240 872 316
rect 888 228 892 332
rect 924 200 928 380
rect 900 196 928 200
rect 932 88 936 203
rect 740 55 744 80
rect 880 52 884 84
rect 996 80 1000 500
rect 1232 404 1236 708
rect 1048 188 1052 276
rect 1072 240 1076 324
rect 1092 228 1096 340
rect 1128 200 1132 388
rect 1232 272 1236 400
rect 1240 336 1244 717
rect 1380 484 1384 621
rect 1676 516 1680 721
rect 1104 196 1132 200
rect 1140 160 1144 203
rect 1120 76 1124 156
rect 920 56 924 76
rect 1120 56 1124 72
rect 1060 52 1080 56
rect 20 -52 24 4
rect 80 -28 84 12
rect 88 -16 92 48
rect -868 -409 -864 -192
rect -724 -329 -720 -232
rect -432 -321 -428 -316
rect -408 -429 -404 -184
rect -356 -397 -352 -200
rect -212 -329 -208 -240
rect 92 -429 96 -172
rect 152 -180 156 4
rect 200 -52 204 4
rect 260 -28 264 12
rect 268 -16 272 48
rect 332 -168 336 4
rect 380 -52 384 4
rect 440 -28 444 12
rect 448 -16 452 48
rect 512 -156 516 4
rect 560 -52 564 4
rect 620 -28 624 12
rect 628 -16 632 48
rect 688 -144 692 4
rect 740 -52 744 4
rect 800 -28 804 12
rect 808 -16 812 48
rect 872 -132 876 4
rect 920 -108 924 8
rect 980 -28 984 12
rect 988 -16 992 48
rect 1012 8 1016 12
rect 1052 -120 1056 4
rect 1140 -52 1144 148
rect 1160 48 1164 256
rect 1228 -16 1232 0
rect 1189 -28 1200 -24
rect 208 -405 212 -208
rect 348 -329 352 -248
rect 652 -429 656 -160
rect 732 -405 736 -216
rect 872 -329 876 -256
rect 592 -433 656 -429
rect 1176 -429 1180 -148
rect 1596 -188 1600 432
rect 1604 -196 1608 424
rect 1612 -204 1616 416
rect 1620 -212 1624 408
rect 1696 404 1700 719
rect 1628 -220 1632 400
rect 1216 -425 1220 -224
rect 1360 -329 1364 -264
rect 1636 -292 1640 400
rect 1696 280 1700 400
rect 1732 344 1736 713
rect 1884 492 1888 620
rect 2188 504 2192 720
rect 1772 352 1776 448
rect 1748 40 1752 284
rect 1652 -429 1656 -136
rect 1772 -228 1776 348
rect 1808 360 1812 456
rect 1784 40 1788 292
rect 1808 -60 1812 356
rect 1844 368 1848 464
rect 1820 40 1824 300
rect 1780 -236 1784 -64
rect 1844 -68 1848 364
rect 1880 376 1884 472
rect 1856 40 1860 308
rect 1788 -244 1792 -72
rect 1880 -76 1884 372
rect 1916 384 1920 480
rect 1892 40 1896 316
rect 1796 -252 1800 -80
rect 1916 -84 1920 380
rect 1952 392 1956 488
rect 1928 40 1932 324
rect 1804 -260 1808 -88
rect 1952 -92 1956 388
rect 2216 48 2220 568
rect 1672 -421 1676 -296
rect 1812 -325 1816 -96
rect 2063 -276 2067 44
rect 2248 -52 2252 788
rect 2264 965 2361 969
rect 2264 552 2268 965
rect 2276 942 2380 946
rect 2276 544 2280 942
rect 2288 904 2412 908
rect 2288 536 2292 904
rect 2300 707 2380 711
rect 2300 528 2304 707
rect 2312 678 2412 682
rect 2312 516 2316 678
rect 2328 500 2380 504
rect 2392 480 2396 481
rect 2308 476 2396 480
rect 2264 315 2364 318
rect 2376 315 2380 318
rect 2264 314 2368 315
rect 2264 136 2268 314
rect 2360 311 2368 314
rect 2376 311 2384 315
rect 2340 307 2348 311
rect 2380 295 2384 311
rect 2276 291 2380 295
rect 2392 307 2424 311
rect 2276 124 2280 291
rect 2392 283 2396 307
rect 2428 295 2436 299
rect 2352 279 2424 283
rect 2392 274 2396 279
rect 2288 253 2412 257
rect 2288 112 2292 253
rect 2400 249 2408 253
rect 2340 245 2344 249
rect 2432 245 2436 249
rect 2348 229 2428 233
rect 2372 204 2376 229
rect 2340 200 2348 204
rect 2360 200 2380 204
rect 2396 200 2415 204
rect 2428 200 2436 204
rect 2352 188 2388 192
rect 2340 172 2348 176
rect 2384 172 2388 188
rect 2412 184 2415 200
rect 2384 168 2424 172
rect 2408 164 2412 168
rect 2400 160 2408 164
rect 2340 156 2344 160
rect 2432 156 2436 160
rect 2348 140 2428 144
rect 2396 121 2400 140
rect 2396 117 2408 121
rect 2340 113 2344 117
rect 2432 113 2436 117
rect 2348 97 2428 101
rect 1604 -433 1656 -429
rect 2120 -428 2124 -124
rect 1844 -468 1848 -460
rect 2112 -848 2116 -500
rect 2156 -840 2160 -112
rect 2212 -645 2216 -184
rect 2220 -467 2224 -172
rect 2228 -438 2232 -160
rect 2236 -240 2240 -148
rect 2244 -203 2248 -136
rect 2252 -176 2256 -124
rect 2264 -147 2268 72
rect 2276 31 2280 84
rect 2288 60 2292 96
rect 2360 80 2364 97
rect 2376 80 2380 82
rect 2360 76 2368 80
rect 2376 76 2384 80
rect 2340 72 2348 76
rect 2380 60 2384 76
rect 2288 56 2380 60
rect 2392 72 2424 76
rect 2392 48 2396 72
rect 2428 60 2436 64
rect 2352 44 2424 48
rect 2372 38 2376 44
rect 2392 40 2396 44
rect 2276 27 2412 31
rect 2400 23 2408 27
rect 2340 19 2344 23
rect 2432 19 2436 23
rect 2348 3 2428 7
rect 2372 -12 2376 -10
rect 2400 -12 2404 3
rect 2340 -16 2348 -12
rect 2360 -16 2380 -12
rect 2400 -16 2415 -12
rect 2428 -16 2436 -12
rect 2352 -28 2388 -24
rect 2340 -44 2348 -40
rect 2384 -44 2388 -28
rect 2412 -32 2415 -16
rect 2384 -48 2424 -44
rect 2408 -52 2412 -48
rect 2400 -56 2408 -52
rect 2340 -60 2344 -56
rect 2432 -60 2436 -56
rect 2348 -76 2428 -72
rect 2392 -90 2396 -76
rect 2392 -94 2408 -90
rect 2340 -98 2344 -94
rect 2432 -98 2436 -94
rect 2348 -114 2428 -110
rect 2360 -127 2364 -114
rect 2360 -131 2368 -127
rect 2376 -131 2384 -127
rect 2340 -135 2348 -131
rect 2380 -147 2384 -131
rect 2264 -151 2380 -147
rect 2392 -135 2424 -131
rect 2392 -159 2396 -135
rect 2428 -147 2436 -143
rect 2352 -163 2424 -159
rect 2392 -168 2396 -163
rect 2320 -172 2396 -168
rect 2252 -180 2364 -176
rect 2244 -207 2380 -203
rect 2236 -244 2408 -240
rect 2400 -249 2408 -244
rect 2228 -442 2381 -438
rect 2220 -471 2412 -467
rect 2212 -649 2380 -645
rect 2392 -668 2396 -662
rect 2320 -672 2368 -668
rect 2380 -672 2396 -668
rect 2308 -752 2368 -748
rect 2376 -752 2380 -736
rect 2376 -840 2380 -816
<< metal2 >>
rect 2252 980 2440 984
rect 2436 962 2440 980
rect 2080 788 2248 792
rect -457 721 -400 725
rect 55 721 116 725
rect 1143 721 1192 725
rect 1627 721 1652 725
rect 2131 720 2188 724
rect 1203 708 1232 712
rect 2156 568 2216 572
rect 2220 568 2340 572
rect -396 548 20 552
rect 24 548 2264 552
rect 120 540 236 544
rect 240 540 2276 544
rect 436 532 676 536
rect 680 532 2288 536
rect 596 524 1192 528
rect 1196 524 2300 528
rect 792 512 1676 516
rect 1680 512 2312 516
rect 1000 500 2188 504
rect 2192 500 2324 504
rect 1888 488 1952 492
rect 1384 480 1916 484
rect 900 472 1880 476
rect 376 464 1844 468
rect -188 456 1808 460
rect -700 448 1772 452
rect -888 432 104 436
rect 108 432 1596 436
rect -388 424 300 428
rect 304 424 1604 428
rect 144 416 468 420
rect 472 416 1612 420
rect 652 408 692 412
rect 696 408 1620 412
rect 1236 400 1628 404
rect 1640 400 1696 404
rect 1132 388 1952 392
rect 928 380 1916 384
rect 744 372 1880 376
rect 556 364 1844 368
rect 384 356 1808 360
rect 188 348 1772 352
rect -344 340 344 344
rect 1096 340 1732 344
rect -844 332 148 336
rect 196 332 512 336
rect 892 332 1240 336
rect 696 324 732 328
rect 1076 324 1928 328
rect 872 316 1892 320
rect 676 308 1856 312
rect 496 300 1820 304
rect 328 292 1784 296
rect 132 284 1748 288
rect 1052 276 1696 280
rect 848 268 1232 272
rect 112 256 704 260
rect 708 256 1056 260
rect 1132 256 1160 260
rect 180 203 204 207
rect 376 203 396 207
rect 544 203 564 207
rect 724 203 748 207
rect 920 203 932 207
rect 1124 203 1140 207
rect 1124 156 1140 160
rect 188 148 719 152
rect 729 148 1096 152
rect 160 132 204 136
rect 208 132 2264 136
rect 344 120 396 124
rect 400 120 2276 124
rect 524 108 564 112
rect 568 108 2288 112
rect 704 96 748 100
rect 752 96 2288 100
rect 884 84 932 88
rect 936 84 2276 88
rect 744 80 788 84
rect 204 76 236 80
rect 384 76 432 80
rect 564 76 592 80
rect 924 76 996 80
rect 1124 72 2264 76
rect 172 68 1076 72
rect 1084 52 1120 56
rect 1184 47 1217 48
rect 1183 44 1217 47
rect 1228 44 1741 48
rect 1751 44 1939 48
rect 1943 44 2063 48
rect 2067 44 2216 48
rect 88 32 92 36
rect 268 32 272 36
rect 448 32 452 36
rect 628 32 632 36
rect 808 32 812 36
rect 988 32 992 36
rect 40 -4 44 2
rect 220 -4 224 2
rect 400 -4 404 1
rect 1072 0 1228 4
rect 580 -4 584 0
rect 760 -4 764 0
rect 940 -4 944 0
rect 40 -8 944 -4
rect 1032 -4 1036 0
rect 1032 -8 1208 -4
rect 92 -20 268 -16
rect 272 -20 448 -16
rect 452 -20 628 -16
rect 632 -20 808 -16
rect 812 -20 988 -16
rect 992 -20 1168 -16
rect 84 -32 260 -28
rect 264 -32 440 -28
rect 444 -32 620 -28
rect 624 -32 800 -28
rect 804 -32 980 -28
rect 984 -32 1196 -28
rect 24 -56 200 -52
rect 204 -56 380 -52
rect 384 -56 560 -52
rect 564 -56 740 -52
rect 744 -56 1140 -52
rect 1144 -56 1161 -52
rect 1183 -56 1216 -52
rect 1223 -56 2248 -52
rect 1784 -64 1808 -60
rect 1792 -72 1844 -68
rect 1800 -80 1880 -76
rect 1808 -88 1916 -84
rect 1816 -96 1952 -92
rect 924 -112 2156 -108
rect 1056 -124 2120 -120
rect 2124 -124 2252 -120
rect 876 -136 1652 -132
rect 1656 -136 2244 -132
rect 692 -148 1176 -144
rect 1180 -148 2236 -144
rect 516 -160 652 -156
rect 656 -160 2228 -156
rect 96 -172 332 -168
rect 336 -172 2220 -168
rect -404 -184 152 -180
rect 156 -184 2212 -180
rect -864 -192 1596 -188
rect -352 -200 1604 -196
rect 212 -208 1612 -204
rect 736 -216 1620 -212
rect 1220 -224 1628 -220
rect -720 -232 1772 -228
rect -208 -240 1780 -236
rect 352 -248 1788 -244
rect 876 -256 1796 -252
rect 1364 -264 1804 -260
rect 1640 -296 1672 -292
rect -448 -381 -447 -377
rect 1676 -425 1677 -421
rect 1220 -429 1224 -425
rect -480 -433 -408 -429
rect 32 -433 92 -429
rect 1120 -433 1176 -429
rect 2056 -432 2120 -428
rect 2012 -500 2112 -496
rect 2304 -748 2308 476
rect 2336 311 2340 481
rect 2336 249 2340 307
rect 2436 299 2440 485
rect 2336 204 2340 245
rect 2392 204 2396 270
rect 2436 249 2440 295
rect 2436 204 2440 245
rect 2336 176 2340 200
rect 2336 160 2340 172
rect 2336 117 2340 156
rect 2336 76 2340 113
rect 2336 23 2340 72
rect 2436 160 2440 200
rect 2436 117 2440 156
rect 2436 64 2440 113
rect 2336 -12 2340 19
rect 2372 -6 2376 34
rect 2436 23 2440 60
rect 2336 -40 2340 -16
rect 2336 -56 2340 -44
rect 2336 -94 2340 -60
rect 2336 -131 2340 -98
rect 2316 -668 2320 -172
rect 2336 -187 2340 -135
rect 2436 -12 2440 19
rect 2436 -56 2440 -16
rect 2436 -94 2440 -60
rect 2436 -143 2440 -98
rect 2436 -188 2440 -147
rect 2336 -677 2340 -664
rect 2436 -677 2440 -664
rect 2336 -759 2340 -746
rect 2436 -757 2440 -744
rect 2160 -844 2376 -840
rect 2436 -848 2440 -828
rect 2116 -852 2440 -848
<< ntransistor >>
rect 2424 301 2428 303
rect 2424 286 2428 288
rect 2428 239 2432 241
rect 2424 194 2428 196
rect 2424 182 2428 184
rect 2428 150 2432 152
rect 2428 107 2432 109
rect 2424 66 2428 68
rect 2424 51 2428 53
rect 2428 13 2432 15
rect 2424 -22 2428 -20
rect 2424 -34 2428 -32
rect 2428 -66 2432 -64
rect 2428 -104 2432 -102
rect 2424 -141 2428 -139
rect 2424 -156 2428 -154
<< ptransistor >>
rect 2348 301 2352 303
rect 2348 286 2352 288
rect 2344 239 2348 241
rect 2348 194 2352 196
rect 2348 182 2352 184
rect 2344 150 2348 152
rect 2344 107 2348 109
rect 2348 66 2352 68
rect 2348 51 2352 53
rect 2344 13 2348 15
rect 2348 -22 2352 -20
rect 2348 -34 2352 -32
rect 2344 -66 2348 -64
rect 2344 -104 2348 -102
rect 2348 -141 2352 -139
rect 2348 -156 2352 -154
<< polycontact >>
rect 2364 307 2368 311
rect 2380 291 2384 295
rect 2408 249 2412 253
rect 2356 200 2360 204
rect 2412 180 2416 184
rect 2408 160 2412 164
rect 2408 117 2412 121
rect 2364 72 2368 76
rect 2380 56 2384 60
rect 2408 23 2412 27
rect 2356 -16 2360 -12
rect 2412 -36 2416 -32
rect 2408 -56 2412 -52
rect 2408 -94 2412 -90
rect 2364 -135 2368 -131
rect 2380 -151 2384 -147
<< ndcontact >>
rect 2424 307 2428 311
rect 2424 295 2428 299
rect 2424 279 2428 283
rect 2428 245 2432 249
rect 2428 229 2432 233
rect 2424 200 2428 204
rect 2424 168 2428 172
rect 2428 156 2432 160
rect 2428 140 2432 144
rect 2428 113 2432 117
rect 2428 97 2432 101
rect 2424 72 2428 76
rect 2424 60 2428 64
rect 2424 44 2428 48
rect 2428 19 2432 23
rect 2428 3 2432 7
rect 2424 -16 2428 -12
rect 2424 -48 2428 -44
rect 2428 -60 2432 -56
rect 2428 -76 2432 -72
rect 2428 -98 2432 -94
rect 2428 -114 2432 -110
rect 2424 -135 2428 -131
rect 2424 -147 2428 -143
rect 2424 -163 2428 -159
<< pdcontact >>
rect 2348 307 2352 311
rect 2348 279 2352 283
rect 2344 245 2348 249
rect 2344 229 2348 233
rect 2348 200 2352 204
rect 2348 188 2352 192
rect 2348 172 2352 176
rect 2344 156 2348 160
rect 2344 140 2348 144
rect 2344 113 2348 117
rect 2344 97 2348 101
rect 2348 72 2352 76
rect 2348 44 2352 48
rect 2344 19 2348 23
rect 2344 3 2348 7
rect 2348 -16 2352 -12
rect 2348 -28 2352 -24
rect 2348 -44 2352 -40
rect 2344 -60 2348 -56
rect 2344 -76 2348 -72
rect 2344 -98 2348 -94
rect 2344 -114 2348 -110
rect 2348 -135 2352 -131
rect 2348 -163 2352 -159
<< m2contact >>
rect 2248 980 2252 984
rect 2248 788 2252 792
rect -400 721 -396 725
rect -892 432 -888 436
rect -848 693 -844 697
rect 116 721 120 725
rect 611 721 615 725
rect -400 548 -396 552
rect -704 448 -700 452
rect -392 424 -388 428
rect -348 689 -344 693
rect -192 456 -188 460
rect 20 548 24 552
rect -348 340 -344 344
rect -848 332 -844 336
rect 116 540 120 544
rect 104 432 108 436
rect 140 416 144 420
rect 192 697 196 701
rect 184 348 188 352
rect 148 332 152 336
rect 128 284 132 288
rect 176 203 180 207
rect 192 332 196 336
rect 236 540 240 544
rect 204 203 208 207
rect 156 132 160 136
rect 204 132 208 136
rect 1192 721 1196 725
rect 1652 721 1656 725
rect 372 464 376 468
rect 432 532 436 536
rect 676 532 680 536
rect 300 424 304 428
rect 380 356 384 360
rect 344 340 348 344
rect 324 292 328 296
rect 372 203 376 207
rect 396 203 400 207
rect 200 76 204 80
rect 236 76 240 80
rect 340 120 344 124
rect 396 120 400 124
rect 592 524 596 528
rect 468 416 472 420
rect 552 364 556 368
rect 512 332 516 336
rect 492 300 496 304
rect 540 203 544 207
rect 564 203 568 207
rect 380 76 384 80
rect 432 76 436 80
rect 520 108 524 112
rect 564 108 568 112
rect 648 408 652 412
rect 692 408 696 412
rect 732 697 736 701
rect 788 512 792 516
rect 692 324 696 328
rect 732 324 736 328
rect 740 372 744 376
rect 672 308 676 312
rect 720 203 724 207
rect 748 203 752 207
rect 560 76 564 80
rect 592 76 596 80
rect 700 96 704 100
rect 748 96 752 100
rect 1240 717 1244 721
rect 1199 708 1203 712
rect 1232 708 1236 712
rect 1192 524 1196 528
rect 896 472 900 476
rect 996 500 1000 504
rect 924 380 928 384
rect 888 332 892 336
rect 868 316 872 320
rect 844 268 848 272
rect 916 203 920 207
rect 932 203 936 207
rect 740 80 744 84
rect 788 80 792 84
rect 880 84 884 88
rect 932 84 936 88
rect 1232 400 1236 404
rect 1128 388 1132 392
rect 1092 340 1096 344
rect 1072 324 1076 328
rect 1048 276 1052 280
rect 1120 203 1124 207
rect 2188 720 2192 724
rect 1676 512 1680 516
rect 1380 480 1384 484
rect 1240 332 1244 336
rect 1596 432 1600 436
rect 1232 268 1236 272
rect 1160 256 1164 260
rect 1140 203 1144 207
rect 920 76 924 80
rect 996 76 1000 80
rect 1120 156 1124 160
rect 1140 156 1144 160
rect 1120 72 1124 76
rect 1080 52 1084 56
rect 1120 52 1124 56
rect 1140 148 1144 152
rect 88 48 92 52
rect 268 48 272 52
rect 88 -20 92 -16
rect 80 -32 84 -28
rect 20 -56 24 -52
rect 92 -172 96 -168
rect -408 -184 -404 -180
rect -868 -192 -864 -188
rect -724 -232 -720 -228
rect -868 -413 -864 -409
rect -356 -200 -352 -196
rect -212 -240 -208 -236
rect -356 -401 -352 -397
rect -408 -433 -404 -429
rect 448 48 452 52
rect 268 -20 272 -16
rect 260 -32 264 -28
rect 200 -56 204 -52
rect 628 48 632 52
rect 448 -20 452 -16
rect 440 -32 444 -28
rect 380 -56 384 -52
rect 808 48 812 52
rect 628 -20 632 -16
rect 620 -32 624 -28
rect 560 -56 564 -52
rect 988 48 992 52
rect 808 -20 812 -16
rect 800 -32 804 -28
rect 740 -56 744 -52
rect 988 -20 992 -16
rect 980 -32 984 -28
rect 920 -112 924 -108
rect 1160 44 1164 48
rect 1228 0 1232 4
rect 1208 -8 1212 -4
rect 1168 -20 1172 -16
rect 1196 -32 1200 -28
rect 1140 -56 1144 -52
rect 1052 -124 1056 -120
rect 872 -136 876 -132
rect 688 -148 692 -144
rect 1176 -148 1180 -144
rect 512 -160 516 -156
rect 652 -160 656 -156
rect 332 -172 336 -168
rect 152 -184 156 -180
rect 208 -208 212 -204
rect 348 -248 352 -244
rect 208 -409 212 -405
rect 732 -216 736 -212
rect 872 -256 876 -252
rect 732 -409 736 -405
rect 92 -433 96 -429
rect 588 -433 592 -429
rect 1596 -192 1600 -188
rect 1604 424 1608 428
rect 1604 -200 1608 -196
rect 1612 416 1616 420
rect 1612 -208 1616 -204
rect 1620 408 1624 412
rect 1620 -216 1624 -212
rect 1628 400 1632 404
rect 1216 -224 1220 -220
rect 1628 -224 1632 -220
rect 1636 400 1640 404
rect 1360 -264 1364 -260
rect 1696 400 1700 404
rect 1732 713 1736 717
rect 2188 500 2192 504
rect 2216 568 2220 572
rect 1884 488 1888 492
rect 1952 488 1956 492
rect 1916 480 1920 484
rect 1880 472 1884 476
rect 1844 464 1848 468
rect 1808 456 1812 460
rect 1732 340 1736 344
rect 1772 448 1776 452
rect 1772 348 1776 352
rect 1696 276 1700 280
rect 1748 284 1752 288
rect 1636 -296 1640 -292
rect 1652 -136 1656 -132
rect 1216 -429 1220 -425
rect 1808 356 1812 360
rect 1784 292 1788 296
rect 1844 364 1848 368
rect 1820 300 1824 304
rect 1772 -232 1776 -228
rect 1780 -64 1784 -60
rect 1808 -64 1812 -60
rect 1880 372 1884 376
rect 1856 308 1860 312
rect 1780 -240 1784 -236
rect 1788 -72 1792 -68
rect 1844 -72 1848 -68
rect 1916 380 1920 384
rect 1892 316 1896 320
rect 1788 -248 1792 -244
rect 1796 -80 1800 -76
rect 1880 -80 1884 -76
rect 1952 388 1956 392
rect 1928 324 1932 328
rect 1796 -256 1800 -252
rect 1804 -88 1808 -84
rect 1916 -88 1920 -84
rect 1804 -264 1808 -260
rect 1812 -96 1816 -92
rect 1952 -96 1956 -92
rect 2063 44 2067 48
rect 2216 44 2220 48
rect 1672 -296 1676 -292
rect 2264 548 2268 552
rect 2276 540 2280 544
rect 2288 532 2292 536
rect 2300 524 2304 528
rect 2312 512 2316 516
rect 2324 500 2328 504
rect 2304 476 2308 480
rect 2336 307 2340 311
rect 2264 132 2268 136
rect 2436 295 2440 299
rect 2392 270 2396 274
rect 2276 120 2280 124
rect 2336 245 2340 249
rect 2436 245 2440 249
rect 2336 200 2340 204
rect 2392 200 2396 204
rect 2436 200 2440 204
rect 2336 172 2340 176
rect 2336 156 2340 160
rect 2436 156 2440 160
rect 2336 113 2340 117
rect 2436 113 2440 117
rect 2288 108 2292 112
rect 2288 96 2292 100
rect 2276 84 2280 88
rect 2248 -56 2252 -52
rect 2264 72 2268 76
rect 2156 -112 2160 -108
rect 2120 -124 2124 -120
rect 1672 -425 1676 -421
rect 1176 -433 1180 -429
rect 1600 -433 1604 -429
rect 2120 -432 2124 -428
rect 2112 -500 2116 -496
rect 2252 -124 2256 -120
rect 2244 -136 2248 -132
rect 2236 -148 2240 -144
rect 2228 -160 2232 -156
rect 2220 -172 2224 -168
rect 2212 -184 2216 -180
rect 2336 72 2340 76
rect 2436 60 2440 64
rect 2372 34 2376 38
rect 2336 19 2340 23
rect 2436 19 2440 23
rect 2372 -10 2376 -6
rect 2336 -16 2340 -12
rect 2436 -16 2440 -12
rect 2336 -44 2340 -40
rect 2336 -60 2340 -56
rect 2436 -60 2440 -56
rect 2336 -98 2340 -94
rect 2436 -98 2440 -94
rect 2336 -135 2340 -131
rect 2436 -147 2440 -143
rect 2316 -172 2320 -168
rect 2316 -672 2320 -668
rect 2304 -752 2308 -748
rect 2156 -844 2160 -840
rect 2376 -844 2380 -840
rect 2112 -852 2116 -848
use CRA6B  CRA6B_0
timestamp 1667778434
transform 1 0 1588 0 1 -509
box -2452 -32 516 241
use CRS6B  CRS6B_0
timestamp 1667778937
transform 1 0 1611 0 -1 801
box -2492 -32 564 241
use ZeroDetection  ZeroDetection_0
timestamp 1665170909
transform 0 -1 2440 -1 0 965
box -4 0 485 104
use ZeroDetection  ZeroDetection_1
timestamp 1665170909
transform 0 -1 2440 -1 0 -184
box -4 0 485 104
use not  not_0
timestamp 1663614877
transform -1 0 1924 0 1 -56
box 8 0 40 104
use not  not_1
timestamp 1663614877
transform -1 0 1960 0 1 -56
box 8 0 40 104
use not  not_2
timestamp 1663614877
transform -1 0 1888 0 1 -56
box 8 0 40 104
use not  not_3
timestamp 1663614877
transform -1 0 1852 0 1 -56
box 8 0 40 104
use not  not_4
timestamp 1663614877
transform -1 0 1780 0 1 -56
box 8 0 40 104
use not  not_5
timestamp 1663614877
transform -1 0 1816 0 1 -56
box 8 0 40 104
use not  not_6
timestamp 1663614877
transform -1 0 1240 0 1 -56
box 8 0 40 104
use not  not_7
timestamp 1663614877
transform -1 0 1200 0 1 -56
box 8 0 40 104
use or  or_0
timestamp 1663598260
transform 0 -1 2440 -1 0 -672
box 0 0 76 104
use or  or_1
timestamp 1663598260
transform 0 -1 2440 -1 0 -752
box 0 0 76 104
use trans4to1  trans4to1_0
timestamp 1667779387
transform 1 0 56 0 1 8
box -56 -8 120 64
use trans4to1  trans4to1_1
timestamp 1667779387
transform 1 0 236 0 1 8
box -56 -8 120 64
use trans4to1  trans4to1_2
timestamp 1667779387
transform 1 0 416 0 1 8
box -56 -8 120 64
use trans4to1  trans4to1_3
timestamp 1667779387
transform 1 0 596 0 1 8
box -56 -8 120 64
use trans4to1  trans4to1_8
timestamp 1667779387
transform 1 0 776 0 1 8
box -56 -8 120 64
use trans4to1  trans4to1_9
timestamp 1667779387
transform 1 0 956 0 1 8
box -56 -8 120 64
use xor  xor_0
timestamp 1663616262
transform 1 0 680 0 1 156
box -36 -8 63 104
use xor  xor_1
timestamp 1663616262
transform 1 0 500 0 1 156
box -36 -8 63 104
use xor  xor_2
timestamp 1663616262
transform 1 0 332 0 1 156
box -36 -8 63 104
use xor  xor_3
timestamp 1663616262
transform 1 0 136 0 1 156
box -36 -8 63 104
use xor  xor_8
timestamp 1663616262
transform 1 0 876 0 1 156
box -36 -8 63 104
use xor  xor_9
timestamp 1663616262
transform 1 0 1080 0 1 156
box -36 -8 63 104
<< labels >>
rlabel metal1 1845 -466 1845 -466 1 Cin
rlabel metal1 1230 -3 1230 -3 1 s0
rlabel metal1 1198 -27 1198 -27 1 s1
rlabel metal1 1774 -18 1774 -18 1 a5
rlabel metal1 1810 -18 1810 -18 1 a4
rlabel metal1 1846 -18 1846 -18 1 a3
rlabel metal1 1882 -18 1882 -18 1 a2
rlabel metal1 1918 -18 1918 -18 1 a1
rlabel metal1 1954 -18 1954 -18 1 a0
rlabel metal1 1598 -18 1598 -18 1 b5
rlabel metal1 1606 -18 1606 -18 1 b4
rlabel metal1 1614 -18 1614 -18 1 b3
rlabel metal1 1622 -18 1622 -18 1 b2
rlabel metal1 1630 -18 1630 -18 1 b1
rlabel metal1 1638 -18 1638 -18 1 b0
rlabel metal1 -430 -318 -430 -318 1 CoutAdd
rlabel metal1 -408 619 -408 619 1 CoutSub
rlabel metal2 90 34 90 34 1 o5
rlabel metal2 270 34 270 34 1 o4
rlabel metal2 450 34 450 34 1 o3
rlabel metal2 630 34 630 34 1 o2
rlabel metal2 810 34 810 34 1 o1
rlabel metal2 1994 -54 1994 -54 1 gnd
rlabel metal2 1998 46 1998 46 1 vdd
rlabel metal2 990 34 990 34 1 o0
<< end >>
